// Evan Harrington
// CSCI320
// Project 1 
////////////// Add4 module /////////////
module add4 (input [31:0] currPC, output [31:0] PCplus4);
	assign PCplus4 = currPC + 4;
endmodule